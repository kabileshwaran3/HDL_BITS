module top_module(
    output zero
);// Module body starts after semicolon
    zero=1'b0;

endmodule
